`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    10:23:07 05/29/2009 
// Design Name: 
// Module Name:    nBitRegister 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////

module Detect_Memory(clock,address,data);

parameter amount=26*26;

input clock;
input[9:0] address;
reg[7:0] mem[0:amount-1];
output reg[7:0] data;


initial begin

mem[0]=0;
mem[1]=0;
mem[2]=0;
mem[3]=0;
mem[4]=0;
mem[5]=0;
mem[6]=0;
mem[7]=0;
mem[8]=0;
mem[9]=0;
mem[10]=0;
mem[11]=0;
mem[12]=0;
mem[13]=0;
mem[14]=0;
mem[15]=0;
mem[16]=0;
mem[17]=0;
mem[18]=0;
mem[19]=0;
mem[20]=0;
mem[21]=0;
mem[22]=0;
mem[23]=0;
mem[24]=0;
mem[25]=0;
mem[26]=0;
mem[27]=255;
mem[28]=255;
mem[29]=255;
mem[30]=255;
mem[31]=255;
mem[32]=255;
mem[33]=255;
mem[34]=255;
mem[35]=255;
mem[36]=255;
mem[37]=255;
mem[38]=255;
mem[39]=255;
mem[40]=255;
mem[41]=255;
mem[42]=255;
mem[43]=255;
mem[44]=255;
mem[45]=0;
mem[46]=0;
mem[47]=0;
mem[48]=0;
mem[49]=0;
mem[50]=0;
mem[51]=0;
mem[52]=0;
mem[53]=255;
mem[54]=255;
mem[55]=255;
mem[56]=255;
mem[57]=255;
mem[58]=255;
mem[59]=255;
mem[60]=255;
mem[61]=255;
mem[62]=255;
mem[63]=255;
mem[64]=255;
mem[65]=255;
mem[66]=255;
mem[67]=255;
mem[68]=255;
mem[69]=255;
mem[70]=255;
mem[71]=0;
mem[72]=0;
mem[73]=0;
mem[74]=0;
mem[75]=0;
mem[76]=0;
mem[77]=0;
mem[78]=0;
mem[79]=255;
mem[80]=255;
mem[81]=0;
mem[82]=0;
mem[83]=0;
mem[84]=255;
mem[85]=255;
mem[86]=255;
mem[87]=255;
mem[88]=255;
mem[89]=255;
mem[90]=255;
mem[91]=255;
mem[92]=0;
mem[93]=0;
mem[94]=0;
mem[95]=255;
mem[96]=255;
mem[97]=0;
mem[98]=0;
mem[99]=0;
mem[100]=0;
mem[101]=0;
mem[102]=0;
mem[103]=0;
mem[104]=0;
mem[105]=255;
mem[106]=255;
mem[107]=0;
mem[108]=255;
mem[109]=0;
mem[110]=255;
mem[111]=255;
mem[112]=255;
mem[113]=255;
mem[114]=255;
mem[115]=255;
mem[116]=255;
mem[117]=255;
mem[118]=0;
mem[119]=255;
mem[120]=0;
mem[121]=255;
mem[122]=255;
mem[123]=0;
mem[124]=0;
mem[125]=0;
mem[126]=0;
mem[127]=0;
mem[128]=0;
mem[129]=0;
mem[130]=0;
mem[131]=255;
mem[132]=255;
mem[133]=0;
mem[134]=0;
mem[135]=0;
mem[136]=255;
mem[137]=255;
mem[138]=255;
mem[139]=255;
mem[140]=255;
mem[141]=255;
mem[142]=255;
mem[143]=255;
mem[144]=0;
mem[145]=0;
mem[146]=0;
mem[147]=255;
mem[148]=255;
mem[149]=0;
mem[150]=0;
mem[151]=0;
mem[152]=0;
mem[153]=0;
mem[154]=0;
mem[155]=0;
mem[156]=0;
mem[157]=255;
mem[158]=255;
mem[159]=255;
mem[160]=255;
mem[161]=255;
mem[162]=255;
mem[163]=255;
mem[164]=255;
mem[165]=255;
mem[166]=255;
mem[167]=255;
mem[168]=255;
mem[169]=255;
mem[170]=255;
mem[171]=255;
mem[172]=255;
mem[173]=255;
mem[174]=255;
mem[175]=0;
mem[176]=0;
mem[177]=0;
mem[178]=0;
mem[179]=0;
mem[180]=0;
mem[181]=0;
mem[182]=0;
mem[183]=255;
mem[184]=255;
mem[185]=255;
mem[186]=255;
mem[187]=255;
mem[188]=255;
mem[189]=255;
mem[190]=255;
mem[191]=255;
mem[192]=255;
mem[193]=255;
mem[194]=255;
mem[195]=255;
mem[196]=255;
mem[197]=255;
mem[198]=255;
mem[199]=255;
mem[200]=255;
mem[201]=0;
mem[202]=0;
mem[203]=0;
mem[204]=0;
mem[205]=0;
mem[206]=0;
mem[207]=0;
mem[208]=0;
mem[209]=255;
mem[210]=255;
mem[211]=255;
mem[212]=255;
mem[213]=255;
mem[214]=255;
mem[215]=255;
mem[216]=255;
mem[217]=255;
mem[218]=255;
mem[219]=255;
mem[220]=255;
mem[221]=255;
mem[222]=255;
mem[223]=255;
mem[224]=255;
mem[225]=255;
mem[226]=255;
mem[227]=0;
mem[228]=0;
mem[229]=0;
mem[230]=0;
mem[231]=0;
mem[232]=0;
mem[233]=0;
mem[234]=0;
mem[235]=255;
mem[236]=255;
mem[237]=255;
mem[238]=255;
mem[239]=255;
mem[240]=255;
mem[241]=255;
mem[242]=255;
mem[243]=0;
mem[244]=0;
mem[245]=255;
mem[246]=255;
mem[247]=255;
mem[248]=255;
mem[249]=255;
mem[250]=255;
mem[251]=255;
mem[252]=255;
mem[253]=0;
mem[254]=0;
mem[255]=0;
mem[256]=0;
mem[257]=0;
mem[258]=0;
mem[259]=0;
mem[260]=0;
mem[261]=255;
mem[262]=255;
mem[263]=255;
mem[264]=255;
mem[265]=255;
mem[266]=255;
mem[267]=255;
mem[268]=255;
mem[269]=0;
mem[270]=0;
mem[271]=255;
mem[272]=255;
mem[273]=255;
mem[274]=255;
mem[275]=255;
mem[276]=255;
mem[277]=255;
mem[278]=255;
mem[279]=0;
mem[280]=0;
mem[281]=0;
mem[282]=0;
mem[283]=0;
mem[284]=0;
mem[285]=0;
mem[286]=0;
mem[287]=255;
mem[288]=255;
mem[289]=255;
mem[290]=255;
mem[291]=255;
mem[292]=255;
mem[293]=255;
mem[294]=255;
mem[295]=255;
mem[296]=255;
mem[297]=255;
mem[298]=255;
mem[299]=255;
mem[300]=255;
mem[301]=255;
mem[302]=255;
mem[303]=255;
mem[304]=255;
mem[305]=0;
mem[306]=0;
mem[307]=0;
mem[308]=0;
mem[309]=0;
mem[310]=0;
mem[311]=0;
mem[312]=0;
mem[313]=255;
mem[314]=255;
mem[315]=255;
mem[316]=255;
mem[317]=255;
mem[318]=255;
mem[319]=255;
mem[320]=255;
mem[321]=255;
mem[322]=255;
mem[323]=255;
mem[324]=255;
mem[325]=255;
mem[326]=255;
mem[327]=255;
mem[328]=255;
mem[329]=255;
mem[330]=255;
mem[331]=0;
mem[332]=0;
mem[333]=0;
mem[334]=0;
mem[335]=0;
mem[336]=0;
mem[337]=0;
mem[338]=0;
mem[339]=255;
mem[340]=255;
mem[341]=255;
mem[342]=255;
mem[343]=255;
mem[344]=255;
mem[345]=255;
mem[346]=255;
mem[347]=255;
mem[348]=255;
mem[349]=255;
mem[350]=255;
mem[351]=255;
mem[352]=255;
mem[353]=255;
mem[354]=255;
mem[355]=255;
mem[356]=255;
mem[357]=0;
mem[358]=0;
mem[359]=0;
mem[360]=0;
mem[361]=0;
mem[362]=0;
mem[363]=0;
mem[364]=0;
mem[365]=255;
mem[366]=255;
mem[367]=255;
mem[368]=255;
mem[369]=255;
mem[370]=255;
mem[371]=0;
mem[372]=0;
mem[373]=0;
mem[374]=0;
mem[375]=0;
mem[376]=0;
mem[377]=255;
mem[378]=255;
mem[379]=255;
mem[380]=255;
mem[381]=255;
mem[382]=255;
mem[383]=0;
mem[384]=0;
mem[385]=0;
mem[386]=0;
mem[387]=0;
mem[388]=0;
mem[389]=0;
mem[390]=0;
mem[391]=255;
mem[392]=255;
mem[393]=255;
mem[394]=255;
mem[395]=255;
mem[396]=255;
mem[397]=0;
mem[398]=255;
mem[399]=255;
mem[400]=255;
mem[401]=255;
mem[402]=0;
mem[403]=255;
mem[404]=255;
mem[405]=255;
mem[406]=255;
mem[407]=255;
mem[408]=255;
mem[409]=0;
mem[410]=0;
mem[411]=0;
mem[412]=0;
mem[413]=0;
mem[414]=0;
mem[415]=0;
mem[416]=0;
mem[417]=255;
mem[418]=255;
mem[419]=255;
mem[420]=255;
mem[421]=255;
mem[422]=255;
mem[423]=0;
mem[424]=255;
mem[425]=255;
mem[426]=255;
mem[427]=255;
mem[428]=0;
mem[429]=255;
mem[430]=255;
mem[431]=255;
mem[432]=255;
mem[433]=255;
mem[434]=255;
mem[435]=0;
mem[436]=0;
mem[437]=0;
mem[438]=0;
mem[439]=0;
mem[440]=0;
mem[441]=0;
mem[442]=0;
mem[443]=255;
mem[444]=255;
mem[445]=255;
mem[446]=255;
mem[447]=255;
mem[448]=255;
mem[449]=0;
mem[450]=0;
mem[451]=0;
mem[452]=0;
mem[453]=0;
mem[454]=0;
mem[455]=255;
mem[456]=255;
mem[457]=255;
mem[458]=255;
mem[459]=255;
mem[460]=255;
mem[461]=0;
mem[462]=0;
mem[463]=0;
mem[464]=0;
mem[465]=0;
mem[466]=0;
mem[467]=0;
mem[468]=0;
mem[469]=255;
mem[470]=255;
mem[471]=255;
mem[472]=255;
mem[473]=255;
mem[474]=255;
mem[475]=255;
mem[476]=255;
mem[477]=255;
mem[478]=255;
mem[479]=255;
mem[480]=255;
mem[481]=255;
mem[482]=255;
mem[483]=255;
mem[484]=255;
mem[485]=255;
mem[486]=255;
mem[487]=0;
mem[488]=0;
mem[489]=0;
mem[490]=0;
mem[491]=0;
mem[492]=0;
mem[493]=0;
mem[494]=0;
mem[495]=0;
mem[496]=0;
mem[497]=0;
mem[498]=0;
mem[499]=0;
mem[500]=0;
mem[501]=0;
mem[502]=0;
mem[503]=0;
mem[504]=0;
mem[505]=0;
mem[506]=0;
mem[507]=0;
mem[508]=0;
mem[509]=0;
mem[510]=0;
mem[511]=0;
mem[512]=0;
mem[513]=0;
mem[514]=0;
mem[515]=0;
mem[516]=0;
mem[517]=0;
mem[518]=0;
mem[519]=0;
mem[520]=0;
mem[521]=0;
mem[522]=0;
mem[523]=0;
mem[524]=0;
mem[525]=0;
mem[526]=0;
mem[527]=0;
mem[528]=0;
mem[529]=0;
mem[530]=0;
mem[531]=0;
mem[532]=0;
mem[533]=0;
mem[534]=0;
mem[535]=0;
mem[536]=0;
mem[537]=0;
mem[538]=0;
mem[539]=0;
mem[540]=0;
mem[541]=0;
mem[542]=0;
mem[543]=0;
mem[544]=0;
mem[545]=0;
mem[546]=0;
mem[547]=0;
mem[548]=0;
mem[549]=0;
mem[550]=0;
mem[551]=0;
mem[552]=0;
mem[553]=0;
mem[554]=0;
mem[555]=0;
mem[556]=0;
mem[557]=0;
mem[558]=0;
mem[559]=0;
mem[560]=0;
mem[561]=0;
mem[562]=0;
mem[563]=0;
mem[564]=0;
mem[565]=0;
mem[566]=0;
mem[567]=0;
mem[568]=0;
mem[569]=0;
mem[570]=0;
mem[571]=0;
mem[572]=0;
mem[573]=0;
mem[574]=0;
mem[575]=0;
mem[576]=0;
mem[577]=0;
mem[578]=0;
mem[579]=0;
mem[580]=0;
mem[581]=0;
mem[582]=0;
mem[583]=0;
mem[584]=0;
mem[585]=0;
mem[586]=0;
mem[587]=0;
mem[588]=0;
mem[589]=0;
mem[590]=0;
mem[591]=0;
mem[592]=0;
mem[593]=0;
mem[594]=0;
mem[595]=0;
mem[596]=0;
mem[597]=0;
mem[598]=0;
mem[599]=0;
mem[600]=0;
mem[601]=0;
mem[602]=0;
mem[603]=0;
mem[604]=0;
mem[605]=0;
mem[606]=0;
mem[607]=0;
mem[608]=0;
mem[609]=0;
mem[610]=0;
mem[611]=0;
mem[612]=0;
mem[613]=0;
mem[614]=0;
mem[615]=0;
mem[616]=0;
mem[617]=0;
mem[618]=0;
mem[619]=0;
mem[620]=0;
mem[621]=0;
mem[622]=0;
mem[623]=0;
mem[624]=0;
mem[625]=0;
mem[626]=0;
mem[627]=0;
mem[628]=0;
mem[629]=0;
mem[630]=0;
mem[631]=0;
mem[632]=0;
mem[633]=0;
mem[634]=0;
mem[635]=0;
mem[636]=0;
mem[637]=0;
mem[638]=0;
mem[639]=0;
mem[640]=0;
mem[641]=0;
mem[642]=0;
mem[643]=0;
mem[644]=0;
mem[645]=0;
mem[646]=0;
mem[647]=0;
mem[648]=0;
mem[649]=0;
mem[650]=0;
mem[651]=0;
mem[652]=0;
mem[653]=0;
mem[654]=0;
mem[655]=0;
mem[656]=0;
mem[657]=0;
mem[658]=0;
mem[659]=0;
mem[660]=0;
mem[661]=0;
mem[662]=0;
mem[663]=0;
mem[664]=0;
mem[665]=0;
mem[666]=0;
mem[667]=0;
mem[668]=0;
mem[669]=0;
mem[670]=0;
mem[671]=0;
mem[672]=0;
mem[673]=0;
mem[674]=0;
mem[675]=0;

end


always@(posedge clock)begin

	data <= mem[address];

end

endmodule

