module histogram (pixel_in,cnt_address, req, counter_out, clk, rst,done );

input[7:0] pixel_in, cnt_address;
output[7:0] counter_out;
input clk, rst, req, done;

// instantiate a CAM-like structure

// SIGNAL DECLARATIONS
wire			done, rst, clk;
reg done, rst, clk;

wire [7:0]		pixel_in;
reg  [7:0]		pixel_in;		// Current state

reg [7:0] counter [255:0]; //counters
reg [7:0] cnt_address;

// MAIN CODE

// Prepare the histogram


always @(posedge clk) begin
if ( rst && ~done )
begin
	case (pixel_in)
		2'b00000000:counter[0] <= counter[0] + 1;	
		2'b00000001:counter[1] <= counter[1] + 1;
		2'b00000010:counter[2] <= counter[2] + 1;	
		2'b00000011:counter[3] <= counter[3] + 1;
		2'b00000100:counter[4] <= counter[4] + 1;
		2'b00000101:counter[5] <= counter[5] + 1;
		2'b00000110:counter[6] <= counter[6] + 1;
		2'b00000111:counter[7] <= counter[7] + 1;
		2'b00001000:counter[8] <= counter[8] + 1;
		2'b00001001:counter[9] <= counter[9] + 1;
		2'b00001010:counter[10] <= counter[10] + 1;
		2'b00001011:counter[11] <= counter[11] + 1;
		2'b00001100:counter[12] <= counter[12] + 1;
		2'b00001101:counter[13] <= counter[13] + 1;
		2'b00001110:counter[14] <= counter[14] + 1;
		2'b00001111:counter[15] <= counter[15] + 1;
		2'b00010000:counter[16] <= counter[16] + 1;
		2'b00010001:counter[17] <= counter[17] + 1;
		2'b00010010:counter[18] <= counter[18] + 1;
		2'b00010011:counter[19] <= counter[19] + 1;
		2'b00010100:counter[20] <= counter[20] + 1;
		2'b00010101:counter[21] <= counter[21] + 1;
		2'b00010110:counter[22] <= counter[22] + 1;
		2'b00010111:counter[23] <= counter[23] + 1;
		2'b00011000:counter[24] <= counter[24] + 1;
		2'b00011001:counter[25] <= counter[25] + 1;
		2'b00011010:counter[26] <= counter[26] + 1;
		2'b00011011:counter[27] <= counter[27] + 1;
		2'b00011100:counter[28] <= counter[28] + 1;
		2'b00011101:counter[29] <= counter[29] + 1;
		2'b00011110:counter[30] <= counter[30] + 1;
		2'b00011111:counter[31] <= counter[31] + 1;
		2'b00100000:counter[32] <= counter[32] + 1;
		2'b00100001:counter[33] <= counter[33] + 1;
		2'b00100010:counter[34] <= counter[34] + 1;
		2'b00100011:counter[35] <= counter[35] + 1;
		2'b00100100:counter[36] <= counter[36] + 1;
		2'b00100101:counter[37] <= counter[37] + 1;
		2'b00100110:counter[38] <= counter[38] + 1;
		2'b00100111:counter[39] <= counter[39] + 1;
		2'b00101000:counter[40] <= counter[40] + 1;
		2'b00101001:counter[41] <= counter[41] + 1;
		2'b00101010:counter[42] <= counter[42] + 1;
		2'b00101011:counter[43] <= counter[43] + 1;
		2'b00101100:counter[44] <= counter[44] + 1;
		2'b00101101:counter[45] <= counter[45] + 1;
		2'b00101110:counter[46] <= counter[46] + 1;
		2'b00101111:counter[47] <= counter[47] + 1;
		2'b00110000:counter[48] <= counter[48] + 1;
		2'b00110001:counter[49] <= counter[49] + 1;
		2'b00110010:counter[50] <= counter[50] + 1;
		2'b00110011:counter[51] <= counter[51] + 1;
		2'b00110100:counter[52] <= counter[52] + 1;
		2'b00110101:counter[53] <= counter[53] + 1;
		2'b00110110:counter[54] <= counter[54] + 1;
		2'b00110111:counter[55] <= counter[55] + 1;
		2'b00111000:counter[56] <= counter[56] + 1;
		2'b00111001:counter[57] <= counter[57] + 1;
		2'b00111010:counter[58] <= counter[58] + 1;
		2'b00111011:counter[59] <= counter[59] + 1;
		2'b00111100:counter[60] <= counter[60] + 1;
		2'b00111101:counter[61] <= counter[61] + 1;
		2'b00111110:counter[62] <= counter[62] + 1;
		2'b00111111:counter[63] <= counter[63] + 1;
		2'b01000000:counter[64] <= counter[64] + 1;
		2'b01000001:counter[65] <= counter[65] + 1;
		2'b01000010:counter[66] <= counter[66] + 1;
		2'b01000011:counter[67] <= counter[67] + 1;
		2'b01000100:counter[68] <= counter[68] + 1;
		2'b01000101:counter[69] <= counter[69] + 1;
		2'b01000110:counter[70] <= counter[70] + 1;
		2'b01000111:counter[71] <= counter[71] + 1;
		2'b01001000:counter[72] <= counter[72] + 1;
		2'b01001001:counter[73] <= counter[73] + 1;
		2'b01001010:counter[74] <= counter[74] + 1;
		2'b01001011:counter[75] <= counter[75] + 1;
		2'b01001100:counter[76] <= counter[76] + 1;
		2'b01001101:counter[77] <= counter[77] + 1;
		2'b01001110:counter[78] <= counter[78] + 1;
		2'b01001111:counter[79] <= counter[79] + 1;
		2'b01010000:counter[80] <= counter[80] + 1;
		2'b01010001:counter[81] <= counter[81] + 1;
		2'b01010010:counter[82] <= counter[82] + 1;
		2'b01010011:counter[83] <= counter[83] + 1;
		2'b01010100:counter[84] <= counter[84] + 1;
		2'b01010101:counter[85] <= counter[85] + 1;
		2'b01010110:counter[86] <= counter[86] + 1;
		2'b01010111:counter[87] <= counter[87] + 1;
		2'b01011000:counter[88] <= counter[88] + 1;
		2'b01011001:counter[89] <= counter[89] + 1;
		2'b01011010:counter[90] <= counter[90] + 1;
		2'b01011011:counter[91] <= counter[91] + 1;
		2'b01011100:counter[92] <= counter[92] + 1;
		2'b01011101:counter[93] <= counter[93] + 1;
		2'b01011110:counter[94] <= counter[94] + 1;
		2'b01011111:counter[95] <= counter[95] + 1;
		2'b01100000:counter[96] <= counter[96] + 1;
		2'b01100001:counter[97] <= counter[97] + 1;
		2'b01100010:counter[98] <= counter[98] + 1;
		2'b01100011:counter[99] <= counter[99] + 1;
		2'b01100100:counter[100] <= counter[100] + 1;
		2'b01100101:counter[101] <= counter[101] + 1;
		2'b01100110:counter[102] <= counter[102] + 1;
		2'b01100111:counter[103] <= counter[103] + 1;
		2'b01101000:counter[104] <= counter[104] + 1;
		2'b01101001:counter[105] <= counter[105] + 1;
		2'b01101010:counter[106] <= counter[106] + 1;
		2'b01101011:counter[107] <= counter[107] + 1;
		2'b01101100:counter[108] <= counter[108] + 1;
		2'b01101101:counter[109] <= counter[109] + 1;
		2'b01101110:counter[110] <= counter[110] + 1;
		2'b01101111:counter[111] <= counter[111] + 1;
		2'b01110000:counter[112] <= counter[112] + 1;
		2'b01110001:counter[113] <= counter[113] + 1;
		2'b01110010:counter[114] <= counter[114] + 1;
		2'b01110011:counter[115] <= counter[115] + 1;
		2'b01110100:counter[116] <= counter[116] + 1;
		2'b01110101:counter[117] <= counter[117] + 1;
		2'b01110110:counter[118] <= counter[118] + 1;
		2'b01110111:counter[119] <= counter[119] + 1;
		2'b01111000:counter[120] <= counter[120] + 1;
		2'b01111001:counter[121] <= counter[121] + 1;
		2'b01111010:counter[122] <= counter[122] + 1;
		2'b01111011:counter[123] <= counter[123] + 1;
		2'b01111100:counter[124] <= counter[124] + 1;
		2'b01111101:counter[125] <= counter[125] + 1;
		2'b01111110:counter[126] <= counter[126] + 1;
		2'b01111111:counter[127] <= counter[127] + 1;
		2'b10000000:counter[128] <= counter[128] + 1;
		2'b10000001:counter[129] <= counter[129] + 1;
		2'b10000010:counter[130] <= counter[130] + 1;
		2'b10000011:counter[131] <= counter[131] + 1;
		2'b10000100:counter[132] <= counter[132] + 1;
		2'b10000101:counter[133] <= counter[133] + 1;
		2'b10000110:counter[134] <= counter[134] + 1;
		2'b10000111:counter[135] <= counter[135] + 1;
		2'b10001000:counter[136] <= counter[136] + 1;
		2'b10001001:counter[137] <= counter[137] + 1;
		2'b10001010:counter[138] <= counter[138] + 1;
		2'b10001011:counter[139] <= counter[139] + 1;
		2'b10001100:counter[140] <= counter[140] + 1;
		2'b10001101:counter[141] <= counter[141] + 1;
		2'b10001110:counter[142] <= counter[142] + 1;
		2'b10001111:counter[143] <= counter[143] + 1;
		2'b10010000:counter[144] <= counter[144] + 1;
		2'b10010001:counter[145] <= counter[145] + 1;
		2'b10010010:counter[146] <= counter[146] + 1;
		2'b10010011:counter[147] <= counter[147] + 1;
		2'b10010100:counter[148] <= counter[148] + 1;
		2'b10010101:counter[149] <= counter[149] + 1;
		2'b10010110:counter[150] <= counter[150] + 1;
		2'b10010111:counter[151] <= counter[151] + 1;
		2'b10011000:counter[152] <= counter[152] + 1;
		2'b10011001:counter[153] <= counter[153] + 1;
		2'b10011010:counter[154] <= counter[154] + 1;
		2'b10011011:counter[155] <= counter[155] + 1;
		2'b10011100:counter[156] <= counter[156] + 1;
		2'b10011101:counter[157] <= counter[157] + 1;
		2'b10011110:counter[158] <= counter[158] + 1;
		2'b10011111:counter[159] <= counter[159] + 1;
		2'b10100000:counter[160] <= counter[160] + 1;
		2'b10100001:counter[161] <= counter[161] + 1;
		2'b10100010:counter[162] <= counter[162] + 1;
		2'b10100011:counter[163] <= counter[163] + 1;
		2'b10100100:counter[164] <= counter[164] + 1;
		2'b10100101:counter[165] <= counter[165] + 1;
		2'b10100110:counter[166] <= counter[166] + 1;
		2'b10100111:counter[167] <= counter[167] + 1;
		2'b10101000:counter[168] <= counter[168] + 1;
		2'b10101001:counter[169] <= counter[169] + 1;
		2'b10101010:counter[170] <= counter[170] + 1;
		2'b10101011:counter[171] <= counter[171] + 1;
		2'b10101100:counter[172] <= counter[172] + 1;
		2'b10101101:counter[173] <= counter[173] + 1;
		2'b10101110:counter[174] <= counter[174] + 1;
		2'b10101111:counter[175] <= counter[175] + 1;
		2'b10110000:counter[176] <= counter[176] + 1;
		2'b10110001:counter[177] <= counter[177] + 1;
		2'b10110010:counter[178] <= counter[178] + 1;
		2'b10110011:counter[179] <= counter[179] + 1;
		2'b10110100:counter[180] <= counter[180] + 1;
		2'b10110101:counter[181] <= counter[181] + 1;
		2'b10110110:counter[182] <= counter[182] + 1;
		2'b10110111:counter[183] <= counter[183] + 1;
		2'b10111000:counter[184] <= counter[184] + 1;
		2'b10111001:counter[185] <= counter[185] + 1;
		2'b10111010:counter[186] <= counter[186] + 1;
		2'b10111011:counter[187] <= counter[187] + 1;
		2'b10111100:counter[188] <= counter[188] + 1;
		2'b10111101:counter[189] <= counter[189] + 1;
		2'b10111110:counter[190] <= counter[190] + 1;
		2'b10111111:counter[191] <= counter[191] + 1;
		2'b11000000:counter[192] <= counter[192] + 1;
		2'b11000001:counter[193] <= counter[193] + 1;
		2'b11000010:counter[194] <= counter[194] + 1;
		2'b11000011:counter[195] <= counter[195] + 1;
		2'b11000100:counter[196] <= counter[196] + 1;
		2'b11000101:counter[197] <= counter[197] + 1;
		2'b11000110:counter[198] <= counter[198] + 1;
		2'b11000111:counter[199] <= counter[199] + 1;
		2'b11001000:counter[200] <= counter[200] + 1;
		2'b11001001:counter[201] <= counter[201] + 1;
		2'b11001010:counter[202] <= counter[202] + 1;
		2'b11001011:counter[203] <= counter[203] + 1;
		2'b11001100:counter[204] <= counter[204] + 1;
		2'b11001101:counter[205] <= counter[205] + 1;
		2'b11001110:counter[206] <= counter[206] + 1;
		2'b11001111:counter[207] <= counter[207] + 1;
		2'b11010000:counter[208] <= counter[208] + 1;
		2'b11010001:counter[209] <= counter[209] + 1;
		2'b11010010:counter[210] <= counter[210] + 1;
		2'b11010011:counter[211] <= counter[211] + 1;
		2'b11010100:counter[212] <= counter[212] + 1;
		2'b11010101:counter[213] <= counter[213] + 1;
		2'b11010110:counter[214] <= counter[214] + 1;
		2'b11010111:counter[215] <= counter[215] + 1;
		2'b11011000:counter[216] <= counter[216] + 1;
		2'b11011001:counter[217] <= counter[217] + 1;
		2'b11011010:counter[218] <= counter[218] + 1;
		2'b11011011:counter[219] <= counter[219] + 1;
		2'b11011100:counter[220] <= counter[220] + 1;
		2'b11011101:counter[221] <= counter[221] + 1;
		2'b11011110:counter[222] <= counter[222] + 1;
		2'b11011111:counter[223] <= counter[223] + 1;
		2'b11100000:counter[224] <= counter[224] + 1;
		2'b11100001:counter[225] <= counter[225] + 1;
		2'b11100010:counter[226] <= counter[226] + 1;
		2'b11100011:counter[227] <= counter[227] + 1;
		2'b11100100:counter[228] <= counter[228] + 1;
		2'b11100101:counter[229] <= counter[229] + 1;
		2'b11100110:counter[230] <= counter[230] + 1;
		2'b11100111:counter[231] <= counter[231] + 1;
		2'b11101000:counter[232] <= counter[232] + 1;
		2'b11101001:counter[233] <= counter[233] + 1;
		2'b11101010:counter[234] <= counter[234] + 1;
		2'b11101011:counter[235] <= counter[235] + 1;
		2'b11101100:counter[236] <= counter[236] + 1;
		2'b11101101:counter[237] <= counter[237] + 1;
		2'b11101110:counter[238] <= counter[238] + 1;
		2'b11101111:counter[239] <= counter[239] + 1;
		2'b11110000:counter[240] <= counter[240] + 1;
		2'b11110001:counter[241] <= counter[241] + 1;
		2'b11110010:counter[242] <= counter[242] + 1;
		2'b11110011:counter[243] <= counter[243] + 1;
		2'b11110100:counter[244] <= counter[244] + 1;
		2'b11110101:counter[245] <= counter[245] + 1;
		2'b11110110:counter[246] <= counter[246] + 1;
		2'b11110111:counter[247] <= counter[247] + 1;
		2'b11111000:counter[248] <= counter[248] + 1;
		2'b11111001:counter[249] <= counter[249] + 1;
		2'b11111010:counter[250] <= counter[250] + 1;
		2'b11111011:counter[251] <= counter[251] + 1;
		2'b11111100:counter[252] <= counter[252] + 1;
		2'b11111101:counter[253] <= counter[253] + 1;
		2'b11111110:counter[254] <= counter[254] + 1;
		2'b11111111:counter[255] <= counter[255] + 1;
		default: newstate <= 8'b00000000;
	endcase
end // end if
else begin
// if done or if reset
counter[0] <= 0;
counter[1] <= 0;
counter[2] <= 0;
counter[3] <= 0;
counter[4] <= 0;
counter[5] <= 0;
counter[6] <= 0;
counter[7] <= 0;
counter[8] <= 0;
counter[9] <= 0;
counter[10] <= 0;
counter[11] <= 0;
counter[12] <= 0;
counter[13] <= 0;
counter[14] <= 0;
counter[15] <= 0;
counter[16] <= 0;
counter[17] <= 0;
counter[18] <= 0;
counter[19] <= 0;
counter[20] <= 0;
counter[21] <= 0;
counter[22] <= 0;
counter[23] <= 0;
counter[24] <= 0;
counter[25] <= 0;
counter[26] <= 0;
counter[27] <= 0;
counter[28] <= 0;
counter[29] <= 0;
counter[30] <= 0;
counter[31] <= 0;
counter[32] <= 0;
counter[33] <= 0;
counter[34] <= 0;
counter[35] <= 0;
counter[36] <= 0;
counter[37] <= 0;
counter[38] <= 0;
counter[39] <= 0;
counter[40] <= 0;
counter[41] <= 0;
counter[42] <= 0;
counter[43] <= 0;
counter[44] <= 0;
counter[45] <= 0;
counter[46] <= 0;
counter[47] <= 0;
counter[48] <= 0;
counter[49] <= 0;
counter[50] <= 0;
counter[51] <= 0;
counter[52] <= 0;
counter[53] <= 0;
counter[54] <= 0;
counter[55] <= 0;
counter[56] <= 0;
counter[57] <= 0;
counter[58] <= 0;
counter[59] <= 0;
counter[60] <= 0;
counter[61] <= 0;
counter[62] <= 0;
counter[63] <= 0;
counter[64] <= 0;
counter[65] <= 0;
counter[66] <= 0;
counter[67] <= 0;
counter[68] <= 0;
counter[69] <= 0;
counter[70] <= 0;
counter[71] <= 0;
counter[72] <= 0;
counter[73] <= 0;
counter[74] <= 0;
counter[75] <= 0;
counter[76] <= 0;
counter[77] <= 0;
counter[78] <= 0;
counter[79] <= 0;
counter[80] <= 0;
counter[81] <= 0;
counter[82] <= 0;
counter[83] <= 0;
counter[84] <= 0;
counter[85] <= 0;
counter[86] <= 0;
counter[87] <= 0;
counter[88] <= 0;
counter[89] <= 0;
counter[90] <= 0;
counter[91] <= 0;
counter[92] <= 0;
counter[93] <= 0;
counter[94] <= 0;
counter[95] <= 0;
counter[96] <= 0;
counter[97] <= 0;
counter[98] <= 0;
counter[99] <= 0;
counter[100] <= 0;
counter[101] <=	0;
counter[102] <=	0;
counter[103] <=	0;
counter[104] <=	0;
counter[105] <=	0;
counter[106] <=	0;
counter[107] <=	0;
counter[108] <=	0;
counter[109] <=	0;
counter[110] <=	0;
counter[111] <=	0;
counter[112] <=	0;
counter[113] <=	0;
counter[114] <=	0;
counter[115] <=	0;
counter[116] <=	0;
counter[117] <=	0;
counter[118] <=	0;
counter[119] <=	0;
counter[120] <=	0;
counter[121] <=	0;
counter[122] <=	0;
counter[123] <=	0;
counter[124] <=	0;
counter[125] <=	0;
counter[126] <=	0;
counter[127] <=	0;
counter[128] <=	0;
counter[129] <=	0;
counter[130] <=	0;
counter[131] <=	0;
counter[132] <=	0;
counter[133] <=	0;
counter[134] <=	0;
counter[135] <=	0;
counter[136] <=	0;
counter[137] <=	0;
counter[138] <=	0;
counter[139] <=	0;
counter[140] <=	0;
counter[141] <=	0;
counter[142] <=	0;
counter[143] <=	0;
counter[144] <=	0;
counter[145] <=	0;
counter[146] <=	0;
counter[147] <=	0;
counter[148] <=	0;
counter[149] <=	0;
counter[150] <=	0;
counter[151] <=	0;
counter[152] <=	0;
counter[153] <=	0;
counter[154] <=	0;
counter[155] <=	0;
counter[156] <=	0;
counter[157] <=	0;
counter[158] <=	0;
counter[159] <=	0;
counter[160] <=	0;
counter[161] <=	0;
counter[162] <=	0;
counter[163] <=	0;
counter[164] <=	0;
counter[165] <=	0;
counter[166] <=	0;
counter[167] <=	0;
counter[168] <=	0;
counter[169] <=	0;
counter[170] <=	0;
counter[171] <=	0;
counter[172] <=	0;
counter[173] <=	0;
counter[174] <=	0;
counter[175] <=	0;
counter[176] <=	0;
counter[177] <=	0;
counter[178] <=	0;
counter[179] <=	0;
counter[180] <=	0;
counter[181] <=	0;
counter[182] <=	0;
counter[183] <=	0;
counter[184] <=	0;
counter[185] <=	0;
counter[186] <=	0;
counter[187] <=	0;
counter[188] <=	0;
counter[189] <=	0;
counter[190] <= 0;
counter[191] <=	0;
counter[192] <=	0;
counter[193] <=	0;
counter[194] <=	0;
counter[195] <=	0;
counter[196] <=	0;
counter[197] <=	0;
counter[198] <=	0;
counter[199] <=	0;
counter[200] <=	0;
counter[201] <=	0;
counter[202] <=	0;
counter[203] <=	0;
counter[204] <=	0;
counter[205] <=	0;
counter[206] <=	0;
counter[207] <=	0;
counter[208] <=	0;
counter[209] <=	0;
counter[210] <=	0;
counter[211] <=	0;
counter[212] <=	0;
counter[213] <=	0;
counter[214] <=	0;
counter[215] <=	0;
counter[216] <=	0;
counter[217] <=	0;
counter[218] <=	0;
counter[219] <=	0;
counter[220] <=	0;
counter[221] <=	0;
counter[222] <=	0;
counter[223] <=	0;
counter[224] <=	0;
counter[225] <=	0;
counter[226] <=	0;
counter[227] <=	0;
counter[228] <=	0;
counter[229] <=	0;
counter[230] <=	0;
counter[231] <=	0;
counter[232] <=	0;
counter[233] <=	0;
counter[234] <=	0;
counter[235] <=	0;
counter[236] <=	0;
counter[237] <=	0;
counter[238] <=	0;
counter[239] <=	0;
counter[240] <=	0;
counter[241] <=	0;
counter[242] <=	0;
counter[243] <=	0;
counter[244] <=	0;
counter[245] <=	0;
counter[246] <=	0;
counter[247] <=	0;
counter[248] <=	0;
counter[249] <=	0;
counter[250] <=	0;
counter[251] <=	0;
counter[252] <=	0;
counter[253] <=	0;
counter[254] <=	0;
counter[255] <=	0;

end // end else

if ( req && done )
begin
counter_out <=counter[cnt_address];
end
else begin
counter_out <=counter_out;
end
  
